`timescale 1p/1ps
/* Horizontal, vertical VGA signals generation
* for 640 x 480 VGA
* */

module HVSync(
    input clk_i,
    input rst_i,
    output hsync_o,
    output vsync_o,
    output display_on,
    output hpos[9:0],
    output vpos[8:0]);




endmodule
