module simpleButton (
    input      button_i,
    output reg led_o
);

assign led_o = button_i;

endmodule
