module simpleButton (
    input      button_i,
    output     led_o
);

assign led_o = button_i;

endmodule
