module servoTop (
    input clk_i,
    output reg srv_o
);

endmodule
